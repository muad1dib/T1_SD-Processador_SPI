// Fazer