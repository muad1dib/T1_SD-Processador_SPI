// Dar uma rechecada nesse negócio


