// Refazer