// Fazer
