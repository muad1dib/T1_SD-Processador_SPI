// Refazer
